configuration na445_circuit_cfg of na445 is
   for circuit
      for all: na444 use configuration work.na444_circuit_cfg;

      end for;
   end for;
end na445_circuit_cfg;

