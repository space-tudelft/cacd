library IEEE;
use IEEE.std_logic_1164.ALL;

entity na447 is
   port(a : in  std_logic;
        b : in  std_logic;
        y : out std_logic);
end na447;

