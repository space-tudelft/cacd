library IEEE;
use IEEE.std_logic_1164.ALL;

PACKAGE param_def IS
constant N : integer;
END param_def;

PACKAGE BODY param_def IS
constant N : integer := 8;
END param_def;

