configuration na444_circuit_cfg of na444 is
   for circuit
   end for;
end na444_circuit_cfg;

