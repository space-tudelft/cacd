library IEEE;
use IEEE.std_logic_1164.ALL;
use WORK.param_def.ALL;

entity na445 is
   port (A:in std_logic;
         B:in std_logic;
         C:in std_logic;
         D:in std_logic;
         Y:out std_logic);
end na445;

