configuration na447_behaviour_cfg of na447 is
   for behaviour
   end for;
end na447_behaviour_cfg;

