

configuration hotel_behaviour_cfg of hotel is
   for behaviour
   end for;
end hotel_behaviour_cfg;


