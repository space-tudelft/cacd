configuration na446_circuit_cfg of na446 is
   for circuit
      for all: na445 use configuration work.na445_circuit_cfg;

      end for;
   end for;
end na446_circuit_cfg;

