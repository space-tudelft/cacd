library IEEE;
use IEEE.std_logic_1164.ALL;


PACKAGE hotel_pkg IS
END hotel_pkg;

