library IEEE;
use IEEE.std_logic_1164.ALL;

entity hotel_tb is
end hotel_tb;
